/home/ise/Desktop/Labratory/PC.vhd